
module reg8 (Latch, CLK, D, Q);
input CLK;
input [7:0] D;
output [7:0] Q;
